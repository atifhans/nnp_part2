// ------------------------------------------//
// Matrix Vector Multiplier Defines Part-1
// ------------------------------------------//
// NAME:  Atif Iqbal
// NETID: aahangar
// SBUID: 111416569
// ------------------------------------------//

package defines_pkg;

    parameter NROWS_A = 3;
    parameter NCOLS_A = 3;
    parameter NROWS_B = 3;
    parameter NCOLS_B = 1;

endpackage
