// ------------------------------------------//
// Matrix Vector Multiplier Defines Part-1
// ------------------------------------------//
// NAME:  Atif Iqbal
// NETID: aahangar
// SBUID: 111416569
// ------------------------------------------//

package defines_pkg;

    parameter NROWS_A = 4;
    parameter NCOLS_A = 4;
    parameter NROWS_B = 4;
    parameter NCOLS_B = 1;

    parameter NUM_S   = 3;
    parameter VEC_S   = 4;

endpackage
